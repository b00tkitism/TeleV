module globals

pub const telegram_api = "https://api.telegram.org/bot"
